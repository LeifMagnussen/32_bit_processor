module AND(A, B, Out);
	input [31:0] A, B;
	output [31:0] Out;
	assign Out = A&B;
endmodule
